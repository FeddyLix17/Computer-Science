module hi(
    input logic[3:0] a
    input logic [1:0] b,
    output logic y
    );
    always_comb
    case (b)
    
endmodule